module main

import os
import term
import args

fn install_packages(global bool) {
    pkg_info := load_package_file()

    println('Installing packages')
    packages := pkg_info.packages

    get_packages(packages, global)
}

fn remove_packages(packages []string) {
    mut removed_packages := []string
    mut lockfile := read_lockfile() or {
        println(err)
        return
    }

    for package in packages {
        pkg_name := if package.starts_with('v-') { package.all_after('v-') } else { package }
        status := delete_package_contents('${ModulesDir}/${pkg_name}')

        if status {
            removed_packages << package
        }
    }

    for package in removed_packages {
        mut pkg_index := 0

        for idx, lock_package in lockfile.packages {
            if lock_package.name == package {
                pkg_index = idx
            }
        }

        lockfile.packages.delete(pkg_index)
    }

    empty_packages := []InstalledPackage

    lockfile.regenerate(empty_packages)

    println('${removed_packages.len} packages were removed.')
}

// TODO: Update packages
fn update_packages() {    
    mut updated_packages := []InstalledPackage

    println('Fetching lockfile')
    mut lockfile := read_lockfile() or {
        println(err)
        create_lockfile()
        return
    }

    println('Updating packages')

    for pkg in lockfile.packages {
        current_hash := pkg.version
        mut latest_hash := current_hash

        os.exec('git --git-dir ${pkg.path}/.git fetch')
        latest_hash = check_git_version(pkg.path)

        if current_hash != latest_hash {
            os.exec('git --git-dir ${pkg.path}/.git pull')

            updated_package := InstalledPackage{
                name: pkg.name,
                path: pkg.path,
                version: latest_hash
            }

            updated_packages << updated_package
        }
    }

    lockfile.regenerate(updated_packages)

    for package in updated_packages {
        println('${package.name}@${package.version}')
    }

    println('${updated_packages.len} packages were updated successfully')
}

fn get_packages(packages []string, global bool) {
    mut installed_packages := []InstalledPackage
    mut lockfile := read_lockfile() or {
        println(err)
        create_lockfile()
        return
    }

    println(lockfile.packages.len)

    for i := 0; i < packages.len; i++ {
        package := get_package(packages[i], global)

        installed_packages << package
    }

    lockfile.regenerate(installed_packages)

    for package in installed_packages {
        println('${package.name}@${package.version}')
    }

    println('${installed_packages.len} packages were installed successfully.')
}

fn show_package_information() {
    pkg_info := load_package_file()
    lockfile := read_lockfile() or {
        println(err)
        create_lockfile()
        return
    }

    dependencies := pkg_info.packages

    println(lockfile.packages.len)

    println('Package name: ${pkg_info.name}')
    println('Dependencies:')
    for i := 0; i < dependencies.len; i++ {
        println('-' + dependencies[i])
    }

    println('\nInstalled packages:\n')

    for i := 0; i < lockfile.packages.len; i++ {
        pkg := lockfile.packages[i]

        println('${pkg.name}')
    }
}

fn show_version() {
    println('vpkg ${Version}')
    println(os.user_os())
}

fn show_help() {
    println('VPkg ${Version}')
    println('An alternative package manager for V.')

    println('\nCOMMANDS\n')

    println('get [packages]                     Fetch and installs packages from the registry or the git repo.')
    println('help                               Prints this help message.')
    println('info                               Show project\'s package information.')
    println('install                            Reads the ".vpkg.json" file and installs the necessary packages.')
    println('remove [packages]                  Removes packages')
    println('update                             Updates packages.')
    println('version                            Prints the Version of this program.')

    println('\nOPTIONS\n')
    println('--global, -g                       Installs the modules/packages into the vlib folder.')
}