// Copyright (c) 2020 vpkg developers
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

module api

import net.urllib

pub interface Provider {
	domains []string
	protocols []string
mut:
	output_dir string
	fetch(url &urllib.URL, folder_name string) ?string
	// get_version returns the version of the package
	get_version(url &urllib.URL) string
	// update updates the package
	update(url &urllib.URL) ?
	// remove removes the package
	remove(url &urllib.URL) ?
}

pub fn (mut pr Provider) set_output_path(output_dir string) {
	pr.output_dir = output_dir
}

pub fn (prs []Provider) find_by_url(url &urllib.URL) ?Provider {
	host := url.host
	scheme := url.scheme

	for _, provider in prs {
		if host in provider.domains || scheme in provider.protocols {
			return provider
		}
	}

	return error('no provider matches the `$scheme` protocol and/or the `$host` domain.')
}